// `default_nettype none
module tt_um_topmodule (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    rca u0 ( // <--- Your module
        .a(a_x),
        .b(b_x),
        .cin(cin_x),
        .sum(sum_x),
        .cout(cout_x)
    );

    // ! DO NOT TOUCH !
    logic [2:0] a_x, b_x, sum_x;
    logic cin_x;
    logic cout_x;

    assign a_x = ui_in[2:0];
    assign b_x = ui_in[5:3];
    assign cin_x = ui_in[6];

    assign uo_out[2:0]  = sum_x;
    assign uo_out[3]    = cout_x;

    assign uo_out[7:4]  = '0;

    assign uio_out      = '0;
    assign uio_oe       = '0;
endmodule
